
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;



entity samirovi_brojaci is
port {
iCLK : in std_logic;
iRESET : std_logic;
iCOUNT : std_logic;
iINC : std_logic;
oCNT1 : std_logic;
oCNT2 : std_logic;
oCMP : std_logic;
end samirovi_brojaci;


architecture Behavioral of samirovi_brojaci is 
 

begin


end Behavioral;

